Library IEEE;
use IEEE.std_logic_1164.all;

entity Bus32to5 is
port (	inputs : in std_logic_vector(31 downto 0);
			s_out : out std_logic_vector(4 downto 0));
end entity;

architecture swag of Bus32to5 is
begin 
	s_out <= 	"00001" when inputs = "00000000000000000000000000000001" else
					"00010" when inputs = "00000000000000000000000000000010" else
					"00011" when inputs = "00000000000000000000000000000100" else
					"00100" when inputs = "00000000000000000000000000001000" else
					"00101" when inputs = "00000000000000000000000000010000" else
					"00110" when inputs = "00000000000000000000000000100000" else
					"00111" when inputs = "00000000000000000000000001000000" else
					"01000" when inputs = "00000000000000000000000010000000" else
					"01001" when inputs = "00000000000000000000000100000000" else
					"01010" when inputs = "00000000000000000000001000000000" else
					"01011" when inputs = "00000000000000000000010000000000" else
					"01100" when inputs = "00000000000000000000100000000000" else
					"01101" when inputs = "00000000000000000001000000000000" else
					"01110" when inputs = "00000000000000000010000000000000" else
					"01111" when inputs = "00000000000000000100000000000000" else
					"10000" when inputs = "00000000000000001000000000000000" else
					"10001" when inputs = "00000000000000010000000000000000" else
					"10010" when inputs = "00000000000000100000000000000000" else
					"10011" when inputs = "00000000000001000000000000000000" else
					"10100" when inputs = "00000000000010000000000000000000" else
					"10101" when inputs = "00000000000100000000000000000000" else
					"10110" when inputs = "00000000001000000000000000000000" else
					"10111" when inputs = "00000000010000000000000000000000" else
					"11000" when inputs = "00000000100000000000000000000000" else
					"00000";
end architecture swag;	


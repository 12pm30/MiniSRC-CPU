-- Copyright (C) 1991-2014 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.4 Build 182 03/12/2014 SJ Web Edition"
-- CREATED		"Mon Feb 15 12:38:10 2016"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY arr_bit_mult IS 
	PORT
	(
		m_in :  IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q_in :  IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		p_out :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END arr_bit_mult;

ARCHITECTURE bdf_type OF arr_bit_mult IS 

COMPONENT arraymultblock
	PORT(PP_in : IN STD_LOGIC;
		 q_in : IN STD_LOGIC;
		 m_in : IN STD_LOGIC;
		 carry_in : IN STD_LOGIC;
		 q_out : OUT STD_LOGIC;
		 carry_out : OUT STD_LOGIC;
		 m_out : OUT STD_LOGIC;
		 PP_Out : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_constant0
	PORT(		 result : OUT STD_LOGIC_VECTOR(0 TO 0)
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_79 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_81 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_85 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_87 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_88 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_89 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_91 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_92 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_95 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_96 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_97 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_98 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_99 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_100 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_101 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_102 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_103 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_104 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_105 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_106 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_107 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_108 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_109 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_110 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_111 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_112 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_113 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_114 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_115 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_116 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_117 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_118 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_119 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_120 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_121 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_122 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_123 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_124 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_125 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_126 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_127 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_128 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_129 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_130 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_131 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_132 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_133 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_134 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_135 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_136 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_137 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_138 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_139 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_140 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_141 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_142 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_143 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_144 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_145 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_146 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_147 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_148 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_149 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_150 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_151 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_152 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_153 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_154 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_155 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_156 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_157 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_158 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_159 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_160 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_161 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_162 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_163 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_164 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_165 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_166 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_167 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_168 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_169 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_170 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_171 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_172 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_173 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_174 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_175 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_176 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_177 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_178 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_179 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_180 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_181 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_182 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_183 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_184 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_185 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_186 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_187 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_188 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_189 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_190 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_191 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_192 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_193 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_194 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_195 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_196 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_197 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_198 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_199 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_200 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_201 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_202 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_203 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_204 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_205 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_206 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_207 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_208 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_209 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_210 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_211 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_212 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_213 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_214 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_215 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_216 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_217 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_218 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_219 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_220 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_221 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_222 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_223 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_224 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_225 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_226 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_227 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_228 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_229 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_230 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_231 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_232 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_233 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_234 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_235 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_236 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_237 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_238 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_239 :  STD_LOGIC;


BEGIN 



b2v_inst : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_0,
		 q_in => SYNTHESIZED_WIRE_1,
		 m_in => m_in(3),
		 carry_in => SYNTHESIZED_WIRE_2,
		 q_out => SYNTHESIZED_WIRE_4,
		 carry_out => SYNTHESIZED_WIRE_5,
		 m_out => SYNTHESIZED_WIRE_12,
		 PP_Out => SYNTHESIZED_WIRE_236);


b2v_inst1 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_3,
		 q_in => SYNTHESIZED_WIRE_4,
		 m_in => m_in(4),
		 carry_in => SYNTHESIZED_WIRE_5,
		 q_out => SYNTHESIZED_WIRE_162,
		 carry_out => SYNTHESIZED_WIRE_163,
		 m_out => SYNTHESIZED_WIRE_124,
		 PP_Out => SYNTHESIZED_WIRE_10);


b2v_inst10 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_6,
		 q_in => SYNTHESIZED_WIRE_7,
		 m_in => SYNTHESIZED_WIRE_8,
		 carry_in => SYNTHESIZED_WIRE_9,
		 q_out => SYNTHESIZED_WIRE_237,
		 carry_out => SYNTHESIZED_WIRE_239,
		 m_out => SYNTHESIZED_WIRE_46,
		 PP_Out => SYNTHESIZED_WIRE_51);


b2v_inst11 : lpm_constant0
PORT MAP(		 result(0) => SYNTHESIZED_WIRE_233);


b2v_inst12 : lpm_constant0
PORT MAP(		 result(0) => SYNTHESIZED_WIRE_86);


b2v_inst13 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_10,
		 q_in => SYNTHESIZED_WIRE_11,
		 m_in => SYNTHESIZED_WIRE_12,
		 carry_in => SYNTHESIZED_WIRE_13,
		 q_out => SYNTHESIZED_WIRE_123,
		 carry_out => SYNTHESIZED_WIRE_125,
		 m_out => SYNTHESIZED_WIRE_34,
		 PP_Out => SYNTHESIZED_WIRE_40);


b2v_inst14 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_14,
		 q_in => q_in(1),
		 m_in => SYNTHESIZED_WIRE_15,
		 carry_in => SYNTHESIZED_WIRE_16,
		 q_out => SYNTHESIZED_WIRE_7,
		 carry_out => SYNTHESIZED_WIRE_9,
		 m_out => SYNTHESIZED_WIRE_52,
		 PP_Out => p_out(1));


b2v_inst15 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_17,
		 q_in => SYNTHESIZED_WIRE_18,
		 m_in => SYNTHESIZED_WIRE_19,
		 carry_in => SYNTHESIZED_WIRE_20,
		 q_out => SYNTHESIZED_WIRE_22,
		 carry_out => SYNTHESIZED_WIRE_24,
		 m_out => SYNTHESIZED_WIRE_56,
		 PP_Out => SYNTHESIZED_WIRE_36);


b2v_inst16 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_21,
		 q_in => SYNTHESIZED_WIRE_22,
		 m_in => SYNTHESIZED_WIRE_23,
		 carry_in => SYNTHESIZED_WIRE_24,
		 q_out => SYNTHESIZED_WIRE_26,
		 carry_out => SYNTHESIZED_WIRE_28,
		 m_out => SYNTHESIZED_WIRE_60,
		 PP_Out => SYNTHESIZED_WIRE_54);


b2v_inst17 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_25,
		 q_in => SYNTHESIZED_WIRE_26,
		 m_in => SYNTHESIZED_WIRE_27,
		 carry_in => SYNTHESIZED_WIRE_28,
		 carry_out => SYNTHESIZED_WIRE_62,
		 m_out => SYNTHESIZED_WIRE_64,
		 PP_Out => SYNTHESIZED_WIRE_58);


b2v_inst18 : lpm_constant0
PORT MAP(		 result(0) => SYNTHESIZED_WIRE_16);


b2v_inst19 : lpm_constant0
PORT MAP(		 result(0) => SYNTHESIZED_WIRE_199);


b2v_inst2 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_29,
		 q_in => SYNTHESIZED_WIRE_30,
		 m_in => m_in(2),
		 carry_in => SYNTHESIZED_WIRE_31,
		 q_out => SYNTHESIZED_WIRE_1,
		 carry_out => SYNTHESIZED_WIRE_2,
		 m_out => SYNTHESIZED_WIRE_238,
		 PP_Out => SYNTHESIZED_WIRE_6);


b2v_inst20 : lpm_constant0
PORT MAP(		 result(0) => SYNTHESIZED_WIRE_161);


b2v_inst21 : lpm_constant0
PORT MAP(		 result(0) => SYNTHESIZED_WIRE_3);


b2v_inst22 : lpm_constant0
PORT MAP(		 result(0) => SYNTHESIZED_WIRE_0);


b2v_inst23 : lpm_constant0
PORT MAP(		 result(0) => SYNTHESIZED_WIRE_29);


b2v_inst24 : lpm_constant0
PORT MAP(		 result(0) => SYNTHESIZED_WIRE_48);


b2v_inst25 : lpm_constant0
PORT MAP(		 result(0) => SYNTHESIZED_WIRE_85);


b2v_inst26 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_32,
		 q_in => SYNTHESIZED_WIRE_33,
		 m_in => SYNTHESIZED_WIRE_34,
		 carry_in => SYNTHESIZED_WIRE_35,
		 q_out => SYNTHESIZED_WIRE_37,
		 carry_out => SYNTHESIZED_WIRE_39,
		 m_out => SYNTHESIZED_WIRE_68,
		 PP_Out => SYNTHESIZED_WIRE_74);


b2v_inst27 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_36,
		 q_in => SYNTHESIZED_WIRE_37,
		 m_in => SYNTHESIZED_WIRE_38,
		 carry_in => SYNTHESIZED_WIRE_39,
		 q_out => SYNTHESIZED_WIRE_55,
		 carry_out => SYNTHESIZED_WIRE_57,
		 m_out => SYNTHESIZED_WIRE_72,
		 PP_Out => SYNTHESIZED_WIRE_66);


b2v_inst28 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_40,
		 q_in => SYNTHESIZED_WIRE_41,
		 m_in => SYNTHESIZED_WIRE_42,
		 carry_in => SYNTHESIZED_WIRE_43,
		 q_out => SYNTHESIZED_WIRE_33,
		 carry_out => SYNTHESIZED_WIRE_35,
		 m_out => SYNTHESIZED_WIRE_76,
		 PP_Out => SYNTHESIZED_WIRE_78);


b2v_inst29 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_44,
		 q_in => SYNTHESIZED_WIRE_45,
		 m_in => SYNTHESIZED_WIRE_46,
		 carry_in => SYNTHESIZED_WIRE_47,
		 q_out => SYNTHESIZED_WIRE_41,
		 carry_out => SYNTHESIZED_WIRE_43,
		 m_out => SYNTHESIZED_WIRE_80,
		 PP_Out => SYNTHESIZED_WIRE_82);


b2v_inst3 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_48,
		 q_in => SYNTHESIZED_WIRE_49,
		 m_in => m_in(1),
		 carry_in => SYNTHESIZED_WIRE_50,
		 q_out => SYNTHESIZED_WIRE_30,
		 carry_out => SYNTHESIZED_WIRE_31,
		 m_out => SYNTHESIZED_WIRE_8,
		 PP_Out => SYNTHESIZED_WIRE_14);


b2v_inst30 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_51,
		 q_in => q_in(2),
		 m_in => SYNTHESIZED_WIRE_52,
		 carry_in => SYNTHESIZED_WIRE_53,
		 q_out => SYNTHESIZED_WIRE_45,
		 carry_out => SYNTHESIZED_WIRE_47,
		 m_out => SYNTHESIZED_WIRE_83,
		 PP_Out => p_out(2));


b2v_inst31 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_54,
		 q_in => SYNTHESIZED_WIRE_55,
		 m_in => SYNTHESIZED_WIRE_56,
		 carry_in => SYNTHESIZED_WIRE_57,
		 q_out => SYNTHESIZED_WIRE_59,
		 carry_out => SYNTHESIZED_WIRE_61,
		 m_out => SYNTHESIZED_WIRE_89,
		 PP_Out => SYNTHESIZED_WIRE_70);


b2v_inst32 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_58,
		 q_in => SYNTHESIZED_WIRE_59,
		 m_in => SYNTHESIZED_WIRE_60,
		 carry_in => SYNTHESIZED_WIRE_61,
		 q_out => SYNTHESIZED_WIRE_63,
		 carry_out => SYNTHESIZED_WIRE_65,
		 m_out => SYNTHESIZED_WIRE_93,
		 PP_Out => SYNTHESIZED_WIRE_87);


b2v_inst33 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_62,
		 q_in => SYNTHESIZED_WIRE_63,
		 m_in => SYNTHESIZED_WIRE_64,
		 carry_in => SYNTHESIZED_WIRE_65,
		 carry_out => SYNTHESIZED_WIRE_95,
		 m_out => SYNTHESIZED_WIRE_97,
		 PP_Out => SYNTHESIZED_WIRE_91);


b2v_inst34 : lpm_constant0
PORT MAP(		 result(0) => SYNTHESIZED_WIRE_53);


b2v_inst35 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_66,
		 q_in => SYNTHESIZED_WIRE_67,
		 m_in => SYNTHESIZED_WIRE_68,
		 carry_in => SYNTHESIZED_WIRE_69,
		 q_out => SYNTHESIZED_WIRE_71,
		 carry_out => SYNTHESIZED_WIRE_73,
		 m_out => SYNTHESIZED_WIRE_101,
		 PP_Out => SYNTHESIZED_WIRE_107);


b2v_inst36 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_70,
		 q_in => SYNTHESIZED_WIRE_71,
		 m_in => SYNTHESIZED_WIRE_72,
		 carry_in => SYNTHESIZED_WIRE_73,
		 q_out => SYNTHESIZED_WIRE_88,
		 carry_out => SYNTHESIZED_WIRE_90,
		 m_out => SYNTHESIZED_WIRE_105,
		 PP_Out => SYNTHESIZED_WIRE_99);


b2v_inst37 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_74,
		 q_in => SYNTHESIZED_WIRE_75,
		 m_in => SYNTHESIZED_WIRE_76,
		 carry_in => SYNTHESIZED_WIRE_77,
		 q_out => SYNTHESIZED_WIRE_67,
		 carry_out => SYNTHESIZED_WIRE_69,
		 m_out => SYNTHESIZED_WIRE_109,
		 PP_Out => SYNTHESIZED_WIRE_111);


b2v_inst38 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_78,
		 q_in => SYNTHESIZED_WIRE_79,
		 m_in => SYNTHESIZED_WIRE_80,
		 carry_in => SYNTHESIZED_WIRE_81,
		 q_out => SYNTHESIZED_WIRE_75,
		 carry_out => SYNTHESIZED_WIRE_77,
		 m_out => SYNTHESIZED_WIRE_113,
		 PP_Out => SYNTHESIZED_WIRE_115);


b2v_inst39 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_82,
		 q_in => q_in(3),
		 m_in => SYNTHESIZED_WIRE_83,
		 carry_in => SYNTHESIZED_WIRE_84,
		 q_out => SYNTHESIZED_WIRE_79,
		 carry_out => SYNTHESIZED_WIRE_81,
		 m_out => SYNTHESIZED_WIRE_116,
		 PP_Out => p_out(3));


b2v_inst4 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_85,
		 q_in => q_in(0),
		 m_in => m_in(0),
		 carry_in => SYNTHESIZED_WIRE_86,
		 q_out => SYNTHESIZED_WIRE_49,
		 carry_out => SYNTHESIZED_WIRE_50,
		 m_out => SYNTHESIZED_WIRE_15,
		 PP_Out => p_out(0));


b2v_inst40 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_87,
		 q_in => SYNTHESIZED_WIRE_88,
		 m_in => SYNTHESIZED_WIRE_89,
		 carry_in => SYNTHESIZED_WIRE_90,
		 q_out => SYNTHESIZED_WIRE_92,
		 carry_out => SYNTHESIZED_WIRE_94,
		 m_out => SYNTHESIZED_WIRE_120,
		 PP_Out => SYNTHESIZED_WIRE_103);


b2v_inst41 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_91,
		 q_in => SYNTHESIZED_WIRE_92,
		 m_in => SYNTHESIZED_WIRE_93,
		 carry_in => SYNTHESIZED_WIRE_94,
		 q_out => SYNTHESIZED_WIRE_96,
		 carry_out => SYNTHESIZED_WIRE_98,
		 m_out => SYNTHESIZED_WIRE_128,
		 PP_Out => SYNTHESIZED_WIRE_118);


b2v_inst42 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_95,
		 q_in => SYNTHESIZED_WIRE_96,
		 m_in => SYNTHESIZED_WIRE_97,
		 carry_in => SYNTHESIZED_WIRE_98,
		 carry_out => SYNTHESIZED_WIRE_130,
		 m_out => SYNTHESIZED_WIRE_132,
		 PP_Out => SYNTHESIZED_WIRE_126);


b2v_inst43 : lpm_constant0
PORT MAP(		 result(0) => SYNTHESIZED_WIRE_84);


b2v_inst44 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_99,
		 q_in => SYNTHESIZED_WIRE_100,
		 m_in => SYNTHESIZED_WIRE_101,
		 carry_in => SYNTHESIZED_WIRE_102,
		 q_out => SYNTHESIZED_WIRE_104,
		 carry_out => SYNTHESIZED_WIRE_106,
		 m_out => SYNTHESIZED_WIRE_136,
		 PP_Out => SYNTHESIZED_WIRE_142);


b2v_inst45 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_103,
		 q_in => SYNTHESIZED_WIRE_104,
		 m_in => SYNTHESIZED_WIRE_105,
		 carry_in => SYNTHESIZED_WIRE_106,
		 q_out => SYNTHESIZED_WIRE_119,
		 carry_out => SYNTHESIZED_WIRE_121,
		 m_out => SYNTHESIZED_WIRE_140,
		 PP_Out => SYNTHESIZED_WIRE_134);


b2v_inst46 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_107,
		 q_in => SYNTHESIZED_WIRE_108,
		 m_in => SYNTHESIZED_WIRE_109,
		 carry_in => SYNTHESIZED_WIRE_110,
		 q_out => SYNTHESIZED_WIRE_100,
		 carry_out => SYNTHESIZED_WIRE_102,
		 m_out => SYNTHESIZED_WIRE_144,
		 PP_Out => SYNTHESIZED_WIRE_146);


b2v_inst47 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_111,
		 q_in => SYNTHESIZED_WIRE_112,
		 m_in => SYNTHESIZED_WIRE_113,
		 carry_in => SYNTHESIZED_WIRE_114,
		 q_out => SYNTHESIZED_WIRE_108,
		 carry_out => SYNTHESIZED_WIRE_110,
		 m_out => SYNTHESIZED_WIRE_148,
		 PP_Out => SYNTHESIZED_WIRE_150);


b2v_inst48 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_115,
		 q_in => q_in(4),
		 m_in => SYNTHESIZED_WIRE_116,
		 carry_in => SYNTHESIZED_WIRE_117,
		 q_out => SYNTHESIZED_WIRE_112,
		 carry_out => SYNTHESIZED_WIRE_114,
		 m_out => SYNTHESIZED_WIRE_151,
		 PP_Out => p_out(4));


b2v_inst49 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_118,
		 q_in => SYNTHESIZED_WIRE_119,
		 m_in => SYNTHESIZED_WIRE_120,
		 carry_in => SYNTHESIZED_WIRE_121,
		 q_out => SYNTHESIZED_WIRE_127,
		 carry_out => SYNTHESIZED_WIRE_129,
		 m_out => SYNTHESIZED_WIRE_155,
		 PP_Out => SYNTHESIZED_WIRE_138);


b2v_inst5 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_122,
		 q_in => SYNTHESIZED_WIRE_123,
		 m_in => SYNTHESIZED_WIRE_124,
		 carry_in => SYNTHESIZED_WIRE_125,
		 q_out => SYNTHESIZED_WIRE_18,
		 carry_out => SYNTHESIZED_WIRE_20,
		 m_out => SYNTHESIZED_WIRE_38,
		 PP_Out => SYNTHESIZED_WIRE_32);


b2v_inst50 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_126,
		 q_in => SYNTHESIZED_WIRE_127,
		 m_in => SYNTHESIZED_WIRE_128,
		 carry_in => SYNTHESIZED_WIRE_129,
		 q_out => SYNTHESIZED_WIRE_131,
		 carry_out => SYNTHESIZED_WIRE_133,
		 m_out => SYNTHESIZED_WIRE_159,
		 PP_Out => SYNTHESIZED_WIRE_153);


b2v_inst51 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_130,
		 q_in => SYNTHESIZED_WIRE_131,
		 m_in => SYNTHESIZED_WIRE_132,
		 carry_in => SYNTHESIZED_WIRE_133,
		 carry_out => SYNTHESIZED_WIRE_164,
		 m_out => SYNTHESIZED_WIRE_166,
		 PP_Out => SYNTHESIZED_WIRE_157);


b2v_inst52 : lpm_constant0
PORT MAP(		 result(0) => SYNTHESIZED_WIRE_117);


b2v_inst53 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_134,
		 q_in => SYNTHESIZED_WIRE_135,
		 m_in => SYNTHESIZED_WIRE_136,
		 carry_in => SYNTHESIZED_WIRE_137,
		 q_out => SYNTHESIZED_WIRE_139,
		 carry_out => SYNTHESIZED_WIRE_141,
		 m_out => SYNTHESIZED_WIRE_170,
		 PP_Out => SYNTHESIZED_WIRE_176);


b2v_inst54 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_138,
		 q_in => SYNTHESIZED_WIRE_139,
		 m_in => SYNTHESIZED_WIRE_140,
		 carry_in => SYNTHESIZED_WIRE_141,
		 q_out => SYNTHESIZED_WIRE_154,
		 carry_out => SYNTHESIZED_WIRE_156,
		 m_out => SYNTHESIZED_WIRE_174,
		 PP_Out => SYNTHESIZED_WIRE_168);


b2v_inst55 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_142,
		 q_in => SYNTHESIZED_WIRE_143,
		 m_in => SYNTHESIZED_WIRE_144,
		 carry_in => SYNTHESIZED_WIRE_145,
		 q_out => SYNTHESIZED_WIRE_135,
		 carry_out => SYNTHESIZED_WIRE_137,
		 m_out => SYNTHESIZED_WIRE_178,
		 PP_Out => SYNTHESIZED_WIRE_180);


b2v_inst56 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_146,
		 q_in => SYNTHESIZED_WIRE_147,
		 m_in => SYNTHESIZED_WIRE_148,
		 carry_in => SYNTHESIZED_WIRE_149,
		 q_out => SYNTHESIZED_WIRE_143,
		 carry_out => SYNTHESIZED_WIRE_145,
		 m_out => SYNTHESIZED_WIRE_182,
		 PP_Out => SYNTHESIZED_WIRE_184);


b2v_inst57 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_150,
		 q_in => q_in(5),
		 m_in => SYNTHESIZED_WIRE_151,
		 carry_in => SYNTHESIZED_WIRE_152,
		 q_out => SYNTHESIZED_WIRE_147,
		 carry_out => SYNTHESIZED_WIRE_149,
		 m_out => SYNTHESIZED_WIRE_185,
		 PP_Out => p_out(5));


b2v_inst58 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_153,
		 q_in => SYNTHESIZED_WIRE_154,
		 m_in => SYNTHESIZED_WIRE_155,
		 carry_in => SYNTHESIZED_WIRE_156,
		 q_out => SYNTHESIZED_WIRE_158,
		 carry_out => SYNTHESIZED_WIRE_160,
		 m_out => SYNTHESIZED_WIRE_189,
		 PP_Out => SYNTHESIZED_WIRE_172);


b2v_inst59 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_157,
		 q_in => SYNTHESIZED_WIRE_158,
		 m_in => SYNTHESIZED_WIRE_159,
		 carry_in => SYNTHESIZED_WIRE_160,
		 q_out => SYNTHESIZED_WIRE_165,
		 carry_out => SYNTHESIZED_WIRE_167,
		 m_out => SYNTHESIZED_WIRE_193,
		 PP_Out => SYNTHESIZED_WIRE_187);


b2v_inst6 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_161,
		 q_in => SYNTHESIZED_WIRE_162,
		 m_in => m_in(5),
		 carry_in => SYNTHESIZED_WIRE_163,
		 q_out => SYNTHESIZED_WIRE_200,
		 carry_out => SYNTHESIZED_WIRE_201,
		 m_out => SYNTHESIZED_WIRE_19,
		 PP_Out => SYNTHESIZED_WIRE_122);


b2v_inst60 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_164,
		 q_in => SYNTHESIZED_WIRE_165,
		 m_in => SYNTHESIZED_WIRE_166,
		 carry_in => SYNTHESIZED_WIRE_167,
		 carry_out => SYNTHESIZED_WIRE_195,
		 m_out => SYNTHESIZED_WIRE_197,
		 PP_Out => SYNTHESIZED_WIRE_191);


b2v_inst61 : lpm_constant0
PORT MAP(		 result(0) => SYNTHESIZED_WIRE_152);


b2v_inst62 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_168,
		 q_in => SYNTHESIZED_WIRE_169,
		 m_in => SYNTHESIZED_WIRE_170,
		 carry_in => SYNTHESIZED_WIRE_171,
		 q_out => SYNTHESIZED_WIRE_173,
		 carry_out => SYNTHESIZED_WIRE_175,
		 m_out => SYNTHESIZED_WIRE_204,
		 PP_Out => SYNTHESIZED_WIRE_210);


b2v_inst63 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_172,
		 q_in => SYNTHESIZED_WIRE_173,
		 m_in => SYNTHESIZED_WIRE_174,
		 carry_in => SYNTHESIZED_WIRE_175,
		 q_out => SYNTHESIZED_WIRE_188,
		 carry_out => SYNTHESIZED_WIRE_190,
		 m_out => SYNTHESIZED_WIRE_208,
		 PP_Out => SYNTHESIZED_WIRE_202);


b2v_inst64 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_176,
		 q_in => SYNTHESIZED_WIRE_177,
		 m_in => SYNTHESIZED_WIRE_178,
		 carry_in => SYNTHESIZED_WIRE_179,
		 q_out => SYNTHESIZED_WIRE_169,
		 carry_out => SYNTHESIZED_WIRE_171,
		 m_out => SYNTHESIZED_WIRE_212,
		 PP_Out => SYNTHESIZED_WIRE_214);


b2v_inst65 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_180,
		 q_in => SYNTHESIZED_WIRE_181,
		 m_in => SYNTHESIZED_WIRE_182,
		 carry_in => SYNTHESIZED_WIRE_183,
		 q_out => SYNTHESIZED_WIRE_177,
		 carry_out => SYNTHESIZED_WIRE_179,
		 m_out => SYNTHESIZED_WIRE_216,
		 PP_Out => SYNTHESIZED_WIRE_218);


b2v_inst66 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_184,
		 q_in => q_in(6),
		 m_in => SYNTHESIZED_WIRE_185,
		 carry_in => SYNTHESIZED_WIRE_186,
		 q_out => SYNTHESIZED_WIRE_181,
		 carry_out => SYNTHESIZED_WIRE_183,
		 m_out => SYNTHESIZED_WIRE_219,
		 PP_Out => p_out(6));


b2v_inst67 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_187,
		 q_in => SYNTHESIZED_WIRE_188,
		 m_in => SYNTHESIZED_WIRE_189,
		 carry_in => SYNTHESIZED_WIRE_190,
		 q_out => SYNTHESIZED_WIRE_192,
		 carry_out => SYNTHESIZED_WIRE_194,
		 m_out => SYNTHESIZED_WIRE_223,
		 PP_Out => SYNTHESIZED_WIRE_206);


b2v_inst68 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_191,
		 q_in => SYNTHESIZED_WIRE_192,
		 m_in => SYNTHESIZED_WIRE_193,
		 carry_in => SYNTHESIZED_WIRE_194,
		 q_out => SYNTHESIZED_WIRE_196,
		 carry_out => SYNTHESIZED_WIRE_198,
		 m_out => SYNTHESIZED_WIRE_227,
		 PP_Out => SYNTHESIZED_WIRE_221);


b2v_inst69 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_195,
		 q_in => SYNTHESIZED_WIRE_196,
		 m_in => SYNTHESIZED_WIRE_197,
		 carry_in => SYNTHESIZED_WIRE_198,
		 carry_out => SYNTHESIZED_WIRE_229,
		 m_out => SYNTHESIZED_WIRE_231,
		 PP_Out => SYNTHESIZED_WIRE_225);


b2v_inst7 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_199,
		 q_in => SYNTHESIZED_WIRE_200,
		 m_in => m_in(6),
		 carry_in => SYNTHESIZED_WIRE_201,
		 q_out => SYNTHESIZED_WIRE_234,
		 carry_out => SYNTHESIZED_WIRE_235,
		 m_out => SYNTHESIZED_WIRE_23,
		 PP_Out => SYNTHESIZED_WIRE_17);


b2v_inst70 : lpm_constant0
PORT MAP(		 result(0) => SYNTHESIZED_WIRE_186);


b2v_inst71 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_202,
		 q_in => SYNTHESIZED_WIRE_203,
		 m_in => SYNTHESIZED_WIRE_204,
		 carry_in => SYNTHESIZED_WIRE_205,
		 q_out => SYNTHESIZED_WIRE_207,
		 carry_out => SYNTHESIZED_WIRE_209,
		 PP_Out => p_out(10));


b2v_inst72 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_206,
		 q_in => SYNTHESIZED_WIRE_207,
		 m_in => SYNTHESIZED_WIRE_208,
		 carry_in => SYNTHESIZED_WIRE_209,
		 q_out => SYNTHESIZED_WIRE_222,
		 carry_out => SYNTHESIZED_WIRE_224,
		 PP_Out => p_out(11));


b2v_inst73 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_210,
		 q_in => SYNTHESIZED_WIRE_211,
		 m_in => SYNTHESIZED_WIRE_212,
		 carry_in => SYNTHESIZED_WIRE_213,
		 q_out => SYNTHESIZED_WIRE_203,
		 carry_out => SYNTHESIZED_WIRE_205,
		 PP_Out => p_out(9));


b2v_inst74 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_214,
		 q_in => SYNTHESIZED_WIRE_215,
		 m_in => SYNTHESIZED_WIRE_216,
		 carry_in => SYNTHESIZED_WIRE_217,
		 q_out => SYNTHESIZED_WIRE_211,
		 carry_out => SYNTHESIZED_WIRE_213,
		 PP_Out => p_out(8));


b2v_inst75 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_218,
		 q_in => q_in(7),
		 m_in => SYNTHESIZED_WIRE_219,
		 carry_in => SYNTHESIZED_WIRE_220,
		 q_out => SYNTHESIZED_WIRE_215,
		 carry_out => SYNTHESIZED_WIRE_217,
		 PP_Out => p_out(7));


b2v_inst76 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_221,
		 q_in => SYNTHESIZED_WIRE_222,
		 m_in => SYNTHESIZED_WIRE_223,
		 carry_in => SYNTHESIZED_WIRE_224,
		 q_out => SYNTHESIZED_WIRE_226,
		 carry_out => SYNTHESIZED_WIRE_228,
		 PP_Out => p_out(12));


b2v_inst77 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_225,
		 q_in => SYNTHESIZED_WIRE_226,
		 m_in => SYNTHESIZED_WIRE_227,
		 carry_in => SYNTHESIZED_WIRE_228,
		 q_out => SYNTHESIZED_WIRE_230,
		 carry_out => SYNTHESIZED_WIRE_232,
		 PP_Out => p_out(13));


b2v_inst78 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_229,
		 q_in => SYNTHESIZED_WIRE_230,
		 m_in => SYNTHESIZED_WIRE_231,
		 carry_in => SYNTHESIZED_WIRE_232,
		 carry_out => p_out(15),
		 PP_Out => p_out(14));


b2v_inst79 : lpm_constant0
PORT MAP(		 result(0) => SYNTHESIZED_WIRE_220);


b2v_inst8 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_233,
		 q_in => SYNTHESIZED_WIRE_234,
		 m_in => m_in(7),
		 carry_in => SYNTHESIZED_WIRE_235,
		 carry_out => SYNTHESIZED_WIRE_25,
		 m_out => SYNTHESIZED_WIRE_27,
		 PP_Out => SYNTHESIZED_WIRE_21);


b2v_inst9 : arraymultblock
PORT MAP(PP_in => SYNTHESIZED_WIRE_236,
		 q_in => SYNTHESIZED_WIRE_237,
		 m_in => SYNTHESIZED_WIRE_238,
		 carry_in => SYNTHESIZED_WIRE_239,
		 q_out => SYNTHESIZED_WIRE_11,
		 carry_out => SYNTHESIZED_WIRE_13,
		 m_out => SYNTHESIZED_WIRE_42,
		 PP_Out => SYNTHESIZED_WIRE_44);


END bdf_type;